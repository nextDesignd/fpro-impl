package env_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import apb_pkg::*;

    // TODO : file name and class name for scoreboard should match
    `include "scoreboard.svh"
    `include "env.svh"
    `include "basic_read_write_seq.svh"

endpackage
