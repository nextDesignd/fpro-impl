`include "apb_if.sv"

package apb_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "apb_txn.svh"
    `include "apb_base_seq.svh"
    `include "apb_slave_driver.svh"
    `include "apb_sequencer.svh"
    `include "apb_master_driver.svh"
    `include "apb_monitor.svh"
    `include "apb_agent.svh"

endpackage

