package env_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import apb_pkg::*;

    `include "env.svh"

endpackage
