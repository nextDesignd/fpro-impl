package env_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import apb_pkg::*;

    `include "env.svh"
    `include "basic_read_write_seq.svh"

endpackage
