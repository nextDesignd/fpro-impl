typedef uvm_sequencer#(apb_txn) apb_sequencer;
